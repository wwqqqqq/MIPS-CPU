`timescale 1ns / 1ps

module top(
input clk,
input [3:0] btn,
input [7:0] sw,
output [3:0] an,
output [7:0] seg,
output [7:0] led
    );


endmodule
