`timescale 1ns / 1ps

module PC(
input clk,
input rst_n,
output pc
    );


endmodule
